




module OLED_ShowData(
	
	input				sys_clk,
	input				rst_n,
	
	
	input				dht11_done,
	input[7:0]	   tempH,	
	input[7:0]	   tempL,
	
    input[7:0]          heart_rate,
    input[7:0]          spo2,           // 【新增】血氧数据
	
	input				ShowData_req,		 //字符显示请求
	input				write_done,			 //iic一组数据写完成
	
	output[23:0]	ShowData_Data,		 //字符显示数据
	
	output			ShowData_finish   //字符显示完成

);


//
//reg[3:0]		tempHH; //tempH的高位
//reg[3:0]		tempHL; //tempH的低位
//reg[3:0]		tempLH;
//reg[3:0]		tempLL;
//
//reg[3:0]		humidityHH;
//reg[3:0]		humidityHL;
//reg[3:0]		humidityLH;
//reg[3:0]		humidityLL;
reg[7:0]        heart_rate_reg;
reg[7:0]        spo2_reg;
reg[7:0]		tempHREG;
reg[7:0]		tempLREG;
reg[7:0]		humidityHREG;
reg[7:0]		humidityLREG;


reg[4:0]	font;

reg[4:0]			font_sel;
reg[4:0] 		font_index;
reg				font_row;

reg[7:0]			show_x;
reg[3:0]			show_y;
reg[23:0]		showfont_data_reg;
wire				onefont_finish;
wire[7:0]		fontdata;

assign onefont_finish  = (font_row == 1'b1 && font_index == 'd10 && write_done == 1'b1) ? 1'b1 : 1'b0;
assign ShowData_finish = (onefont_finish == 1'b1 && font_sel == 'd8) ? 1'b1 : 1'b0;
assign ShowData_Data = showfont_data_reg;

always@(*)
begin
	case(font_index)
	'd0:	showfont_data_reg <= {8'h78,8'h00,8'hB0 + show_y + font_row};
	'd1:  showfont_data_reg <= {8'h78,8'h00,8'h00 + show_x[3:0]};
	'd2:  showfont_data_reg <= {8'h78,8'h00,8'h10 + show_x[7:4]};
	default:	showfont_data_reg <= {8'h78,8'h40,fontdata}; //fontdata
	endcase
end

always@(posedge sys_clk or negedge rst_n)
begin
	if(rst_n == 1'b0)
		font_index <= 'd0;
	else if(write_done == 1'b1 && font_index == 'd10)
		font_index <= 'd0;
	else if(write_done == 1'b1 && ShowData_req == 1'b1)
		font_index <= font_index + 1'b1;
	else
		font_index <= font_index;
end

always@(posedge sys_clk or negedge rst_n)
begin
	if(rst_n == 1'b0)
		font_row <= 1'b0;
	else if(onefont_finish == 1'b1)
		font_row <= 1'b0;
	else if(write_done == 1'b1 && font_index == 'd10)
		font_row <= 1'b1;
	else
		font_row <= font_row;
end


always@(posedge sys_clk or negedge rst_n)
begin
	if(rst_n == 1'b0)
		font_sel <= 'd0;
	else if(ShowData_finish == 1'b1)
		font_sel <= 'd0;
	else if(onefont_finish == 1'b1)
		font_sel <= font_sel + 1'b1;
	else
		font_sel <= font_sel;
end


always@(posedge sys_clk or negedge rst_n)
begin
	if(rst_n == 1'b0)
	begin
		show_x <= 'd0;
		show_y <= 'd0;
	end
    // --- Row 0: 血氧 (font_sel 0,1,2) ---
    else if(font_sel == 'd0) 
	begin 
	    show_x <= 'd54; 
		show_y <= 'd0; 
	end // 百位 (可选)
    else if(font_sel == 'd1) 
	begin 
	    show_x <= 'd62; 
		show_y <= 'd0; 
	end // 十位
    else if(font_sel == 'd2) begin show_x <= 'd70; show_y <= 'd0; end // 个位
    
    // --- Row 3: 温度 (font_sel 3,4,5) ---
    else if(font_sel == 'd3) begin show_x <= 'd54; show_y <= 'd3; end
    else if(font_sel == 'd4) begin show_x <= 'd62; show_y <= 'd3; end
    else if(font_sel == 'd5) begin show_x <= 'd79; show_y <= 'd3; end // 小数
    
    // --- Row 5: 心率 (font_sel 6,7,8) ---
    else if(font_sel == 'd6) begin show_x <= 'd54; show_y <= 'd5; end
    else if(font_sel == 'd7) begin show_x <= 'd62; show_y <= 'd5; end
    else if(font_sel == 'd8) begin show_x <= 'd70; show_y <= 'd5; end
    

	else
	begin
		show_x <= 'd0;
		show_y <= 'd0;
	end
end



always@(posedge sys_clk or negedge rst_n)
begin
	if(rst_n == 1'b0)
		font <= 'd0;
    // 血氧
    else if(font_sel == 'd0) font <= spo2_reg / 100;
    else if(font_sel == 'd1) font <= (spo2_reg / 10) % 10;
    else if(font_sel == 'd2) font <= spo2_reg % 10;
    
    // 温度
    else if(font_sel == 'd3) font <= tempHREG / 10;
    else if(font_sel == 'd4) font <= tempHREG % 10;
    else if(font_sel == 'd5) font <= tempLREG;
    
    // 心率
    else if(font_sel == 'd6) font <= heart_rate_reg / 100;
    else if(font_sel == 'd7) font <= (heart_rate_reg / 10) % 10;
    else if(font_sel == 'd8) font <= heart_rate_reg % 10;
	else
		font <= font;		
end


always@(posedge sys_clk or negedge rst_n)
begin
    if(!rst_n) begin tempHREG<=0; tempLREG<=0; heart_rate_reg<=0; spo2_reg<=0; end
    else if(dht11_done) begin
        tempHREG <= tempH;
        tempLREG <= tempL;
        heart_rate_reg <= heart_rate;
        spo2_reg <= spo2;
    end
end

OLED_NumData OLED_NumDataHP(

	.sys_clk		(sys_clk),
	.rst_n		(rst_n),
	
	.font_row	(font_row),
	.font_sel	(font),
	.index		(font_index - 'd3),
	
	.data			(fontdata)

);

endmodule 